module ysyx_22040759_32add(
    input  [31:0]     a,
    input  [31:0]     b,
    output [31:0]     c
    );
    assign c = a + b;
endmodule
